Example Output
text
[GEN] : Data send to Driver a:4 and b:1
[DRV] : Interface triggered with a:4 and b:1
[MON] : Data send to Scoreboard a:4, b:1 and sum:5
[SCO] : Test Passed for a=4, b=1, sum=5
[ASSERT] SUM_CHECK Pass: Sum:5
🧪 Test Cases
Basic arithmetic operations

Reset functionality verification

Boundary value testing (overflow prevention)

Randomized input testing

Unknown value handling

📈 Verification Metrics
Functional Coverage: 100% for specified constraints

Assertion Coverage: All SVA properties verified

Bug Detection: Catches timing and arithmetic errors

Reset Recovery: Proper reset behavior verified

🎓 Learning Outcomes
This project demonstrates:

Synchronous design principles

Assertion-Based Verification methodology

UVM-style testbench architecture

Constrained random testing

Debugging techniques with SVA

🤝 Contributing
Feel free to:

Add more assertion properties

Extend constraint ranges

Implement functional coverage

Add different adder architectures
